`timescale 1ns / 1ps

module Pipelined_Processor(
    input clk,
    input reset
);

wire [31:0] I1, ALU_Result;
wire [31:0] Instruction_Code, PC, PC1, RD_2, PC_Final, Instruction_Code_1;
reg [31:0] PC_New;
wire [4:0] Rs, Rd, Rt, Write_Reg_Final, wr1, wr2, W1,Rd1, Rs1, Rt1, Rs_New, Rt_New;
wire [31:0] Write_Data_Final, Read_Data_1, Read_Data_2, RD1, RD2, SE1, SE2, A1, Data1, Read_New,
Read_New_1, Data_New_1, Read_FD_Rs, Read_FD_Rt;

wire [31:0] Extended_Offset;
wire Zero, Z1;
wire [15:0] imm;
reg [15:0] Shift;

//Control Unit
wire [5:0] ALU_Op, ALU_Op1;
wire  ALU_Src, Reg_Dest, Is_Branch, Mem_Wr, Mem_Rd, Reg_Wr, Mem_To_Reg;
wire  ALU_Src1, Reg_Dest1, Mem_Wr1, Mem_Rd1, Reg_Wr1, Mem_To_Reg1;
wire  Reg_Dest2, Mem_Wr2, Mem_Rd2, Reg_Wr2, Mem_To_Reg2;
wire  Reg_Wr3, Mem_To_Reg3;

wire [1:0] Forward_Rs, Forward_Rt;

//Stall
wire Stall, clk_Stall;
wire [31:0] I_New;
//----------------------------------------------------------------------------------------
//32-bit instruction code
Instruction_Fetch Fetch1 (clk, reset, Instruction_Code, Is_Branch, PC_New, PC, Stall);

//----------------------------------------------------------------------------------------
//IFD has Instruction_Code as input and Rs,Rt,Rd,immediate data
IFD IFD1(clk,Instruction_Code_1, PC, Rs, Rt, Rd, imm, PC1, I1, Is_Branch);
//Passing same instruction in case of Stall
MUX_Fwd #(31) Instr_1(Instruction_Code, I1, Stall, Instruction_Code_1);

Control_Unit C1(I_New, ALU_Op, ALU_Src, Reg_Dest,
 Is_Branch, Mem_Wr, Mem_Rd, Reg_Wr, Mem_To_Reg);
 
 //To choose Destination Register
 MUX #(4)Dest1 (Rt, Rd, Reg_Dest, Rd1);
 
//Register file
Register_File RFile1 (reset, Rs, Rt, Read_Data_1, Read_Data_2, Write_Reg_Final, Write_Data_Final, Reg_Wr3);
//Sign Extension
Sign_Extend S1 (imm,Extended_Offset);
//Shift left by 2
Shift_Left_2 sl1(Extended_Offset, SE1);

//PC_New value is used for Jump Instruction
always @(PC1, SE1) PC_New = PC1 + SE1;

//----------------------------------------------------------------------------------------
//IDE
IDE IDE1(clk, Read_Data_1, Read_Data_2, Extended_Offset,Rd1, RD1, RD2, SE2,wr1,
ALU_Op, ALU_Src, Reg_Dest, Mem_Wr, Mem_Rd, Reg_Wr, Mem_To_Reg,
ALU_Op1, ALU_Src1, Reg_Dest1, Mem_Wr1, Mem_Rd1, Reg_Wr1, Mem_To_Reg1,
Rs, Rt, Rs1, Rt1);

//Execution Unit
always @(SE2) Shift = SE2[15:0];
//Execution Unit Contains ALU
EXE E1( Read_FD_Rs, Read_FD_Rt, SE2, Shift, wr1, Zero, ALU_Result, RD_2, wr2, ALU_Op1, ALU_Src1);

//----------------------------------------------------------------------------------------
//EXMEM
EXMEM EM1(clk, Zero, ALU_Result, RD_2, wr2, Z1, A1, Data1, W1,
Reg_Dest1, Mem_Wr1, Mem_Rd1, Reg_Wr1, Mem_To_Reg1,
Reg_Dest2, Mem_Wr2, Mem_Rd2, Reg_Wr2, Mem_To_Reg2);

//Data Memory
Data_Memory DM1 (reset, A1, Data1, Read_New, Mem_Rd2, Mem_Wr2);//RD/WR control signal

//----------------------------------------------------------------------------------------
//MEMWB
MEMWB MW1 (clk, Read_New, A1, W1, Read_New_1, Data_New_1, Write_Reg_Final,
Reg_Wr2, Mem_To_Reg2, Reg_Wr3, Mem_To_Reg3);
//TO choose whether there is Memory to Register Transfer
MUX M1 (Data_New_1, Read_New_1, Mem_To_Reg3, Write_Data_Final);

//----------------------------------------------------------------------------------------
//Forwarding Unit
Forward_Unit F1(Rs_New, Rt_New, Reg_Wr2, Reg_Wr3, W1, Write_Reg_Final, Forward_Rs, Forward_Rt);

//Using appropriate data as ALU i/p with usage of Control signals generated by forwarding unit
MUX_2 FD_Rs(RD1, A1, Write_Data_Final, 32'd0, Forward_Rs, Read_FD_Rs);
MUX_2 FD_Rt(RD2, A1, Write_Data_Final, 32'd0, Forward_Rt, Read_FD_Rt);

//In case of stall: Pass Rs=Rt=0, to avoid unnecessary forwarding
MUX_Fwd #(4) Fwd_Stall(Rs1, 5'd0, Stall, Rs_New);
MUX_Fwd #(4) Fwd_Stall1(Rt1, 5'd0, Stall, Rt_New);

//----------------------------------------------------------------------------------------
//Stalling Unit
Stall_Unit Stall_1(Mem_Rd1, Rt1, Rs, Rt, Stall);
//Inserts I_New = 32'd0 so that Control Unit generate all Control Signals as zero
MUX #(31) Instr_stall(I1, 32'd0, Stall, I_New);

endmodule
